CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 120 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 176 457 273
110100498 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 882 108 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5881 0 0
2
43530.4 0
0
2 +V
167 190 268 0 1 3
0 16
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3275 0 0
2
43530.4 1
0
6 74112~
219 648 352 0 7 32
0 16 14 17 14 16 18 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
4203 0 0
2
5.89884e-315 0
0
6 74112~
219 495 351 0 7 32
0 16 15 17 15 16 19 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U4A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
3440 0 0
2
5.89884e-315 5.26354e-315
0
6 74112~
219 333 351 0 7 32
0 16 3 17 3 16 20 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
9102 0 0
2
5.89884e-315 5.30499e-315
0
6 74112~
219 190 351 0 7 32
0 16 16 17 16 16 21 3
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
5586 0 0
2
5.89884e-315 5.32571e-315
0
9 CC 7-Seg~
183 801 141 0 17 19
10 4 5 6 7 8 9 10 22 2
1 1 1 1 0 0 1 2
0
0 0 21088 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
525 0 0
2
5.89884e-315 5.34643e-315
0
6 74LS48
188 802 331 0 14 29
0 13 12 11 3 23 24 10 9 8
7 6 5 4 25
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
6206 0 0
2
5.89884e-315 5.3568e-315
0
9 2-In AND~
219 581 186 0 3 22
0 15 12 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3418 0 0
2
5.89884e-315 5.36716e-315
0
9 2-In AND~
219 420 177 0 3 22
0 3 11 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9312 0 0
2
5.89884e-315 5.37752e-315
0
7 Pulser~
4 65 333 0 10 12
0 26 27 28 17 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7419 0 0
2
5.89884e-315 5.38788e-315
0
37
9 1 2 0 0 4240 0 7 1 0 0 3
801 99
882 99
882 102
0 1 3 0 0 8192 0 0 10 3 0 4
268 316
269 316
269 168
396 168
4 0 3 0 0 0 0 5 0 0 30 3
309 333
268 333
268 315
13 1 4 0 0 8320 0 8 7 0 0 5
834 349
903 349
903 189
780 189
780 177
12 2 5 0 0 8320 0 8 7 0 0 5
834 340
893 340
893 199
786 199
786 177
11 3 6 0 0 8320 0 8 7 0 0 5
834 331
884 331
884 210
792 210
792 177
10 4 7 0 0 8320 0 8 7 0 0 5
834 322
875 322
875 220
798 220
798 177
9 5 8 0 0 8320 0 8 7 0 0 5
834 313
865 313
865 231
804 231
804 177
8 6 9 0 0 16512 0 8 7 0 0 5
834 304
856 304
856 242
810 242
810 177
7 7 10 0 0 16512 0 8 7 0 0 5
834 295
847 295
847 252
816 252
816 177
0 4 3 0 0 8320 0 0 8 30 0 5
225 315
225 477
755 477
755 322
770 322
0 3 11 0 0 8320 0 0 8 24 0 5
368 315
368 469
747 469
747 313
770 313
0 2 12 0 0 8320 0 0 8 22 0 5
531 315
531 460
738 460
738 304
770 304
0 1 13 0 0 12416 0 0 8 29 0 5
685 316
685 452
729 452
729 295
770 295
2 0 14 0 0 4096 0 3 0 0 16 2
624 316
612 316
4 3 14 0 0 8320 0 3 9 0 0 4
624 334
612 334
612 186
602 186
2 0 15 0 0 4096 0 4 0 0 18 2
471 315
458 315
4 0 15 0 0 8320 0 4 0 0 23 3
471 333
458 333
458 177
2 0 16 0 0 4096 0 6 0 0 20 2
166 315
153 315
4 1 16 0 0 8192 0 6 2 0 0 4
166 333
153 333
153 277
190 277
0 0 16 0 0 4096 0 0 0 27 37 2
244 277
244 387
2 7 12 0 0 0 0 9 4 0 0 4
557 195
540 195
540 315
519 315
3 1 15 0 0 0 0 10 9 0 0 2
441 177
557 177
2 7 11 0 0 0 0 10 5 0 0 3
396 186
396 315
357 315
1 0 16 0 0 0 0 5 0 0 27 2
333 288
333 277
1 0 16 0 0 0 0 4 0 0 27 2
495 288
495 277
1 1 16 0 0 4224 0 2 3 0 0 3
190 277
648 277
648 289
1 1 16 0 0 0 0 2 6 0 0 2
190 277
190 288
7 0 13 0 0 0 0 3 0 0 0 2
672 316
711 316
7 2 3 0 0 0 0 6 5 0 0 2
214 315
309 315
3 0 17 0 0 8192 0 4 0 0 34 3
465 324
451 324
451 414
3 0 17 0 0 0 0 5 0 0 34 3
303 324
288 324
288 414
3 0 17 0 0 0 0 6 0 0 34 3
160 324
145 324
145 414
4 3 17 0 0 12416 0 11 3 0 0 6
95 333
117 333
117 414
603 414
603 325
618 325
5 0 16 0 0 0 0 4 0 0 37 2
495 363
495 387
5 0 16 0 0 0 0 5 0 0 37 2
333 363
333 387
5 5 16 0 0 0 0 6 3 0 0 4
190 363
190 387
648 387
648 364
3
-16 0 0 0 400 0 0 0 0 3 2 1 18
7 Georgia
0 0 0 9
9 37 105 64
19 45 94 64
9 BSCPE 1-B
-19 0 0 0 400 0 0 0 0 3 2 1 18
7 Georgia
0 0 0 35
270 56 677 89
280 64 666 87
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
-16 0 0 0 400 0 0 0 0 3 2 1 18
7 Georgia
0 0 0 24
9 11 239 38
19 18 228 37
24 RAMIREZ, MARIA FLIONA A.
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
